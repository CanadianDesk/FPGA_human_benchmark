
//TOP LEVEL MODULE FOR VGA ENCODER

//NEEDS INPUTS:
////1: 2 bits, 00 if Menu, 01 of React, 10 if Chimp, 11 if somethings fucked up 


module zVGAencoder (

);

endmodule   