module VGAreaction();


endmodule