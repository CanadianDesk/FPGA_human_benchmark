module topLevel ();
    
endmodule

