

//TOP LEVEL MODULE FOR VGA ENCODER

//NEEDS INPUTS:
//1) From mainMenu a 2 bit in put based on what is being displayed 0-menu, 1-react, 2-chimp


module zVGAencoder (
    ports
);
    
endmodule