module VGAmenu(
    input clk,
    input iEnable,
    output oEnable,
);



endmodule;