module VGAmenu();



endmodule;