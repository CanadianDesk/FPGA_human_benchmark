



// INPUTS: Reset, clk, mouseX, mouseY
// OUTPUTS: BoxX, BoxY

module (input iReset, clk, [9:0] mouseX, [8:0] mouseY, output [2:0] BoxX, [2:0] BoxY);

endmodule