// Main Menu Key
// Jonah Diamond
// ECE241 Project

// INPUTS
//// 1. 1 bit, whether KEY[0] is pressed
// OUTPUTS
//// idk tbh

// module key0DE1SOC(input KEY[0]);
//     mainMenu mM(.iKey0(KEY[0]));
//     chimp c1(.iKey0(KEY[0]));
// endmodule