//FSM THAT CONTROLS THE VGA


module VGAcontrol();



endmodule;

