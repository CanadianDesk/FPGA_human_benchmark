module mainMenuDataPath();

endmodule